module main
    ( input [7:0] data
    , input spi_clk
    , input mosi
    , output miso
    );

endmodule
